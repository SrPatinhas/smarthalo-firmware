** Profile: "DummyLoad2A_TB-DCSweepVRef"  [ C:\Users\sgelinas\Documents\Git SmartHalo\Hardware\Simulation\electronicload-pspicefiles\dummyload2a_tb\dcsweepvref.sim ] 

** Creating circuit file "DCSweepVRef.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../electronicload-pspicefiles/electronicload.lib" 
* From [PSPICE NETLIST] section of C:\Users\sgelinas\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM VREF 0Vdc 5Vdc 0.1Vdc 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\DummyLoad2A_TB.net" 


.END
