** Profile: "CENTRALLED_TB-trans"  [ C:\Users\sgelinas\Documents\Git SmartHalo\Hardware\Simulation\CentralLEDDriver-PSpiceFiles\CENTRALLED_TB\trans.sim ] 

** Creating circuit file "trans.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../centralleddriver-pspicefiles/centralleddriver.lib" 
* From [PSPICE NETLIST] section of C:\Users\sgelinas\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 10u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\CENTRALLED_TB.net" 


.END
