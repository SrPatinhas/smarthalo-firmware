** Profile: "BATMON_TB-ILOADSWEEP"  [ C:\Users\sgelinas\Documents\Git SmartHalo\Hardware\Simulation\batmon-pspicefiles\batmon_tb\iloadsweep.sim ] 

** Creating circuit file "ILOADSWEEP.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\sgelinas\cdssetup\OrCAD_PSpice/16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN PARAM ILOAD -1.0Adc 1.5Adc 0.25 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\BATMON_TB.net" 


.END
